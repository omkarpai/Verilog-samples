module stimulus_rcfa4
reg [3:0] a,b;